library verilog;
use verilog.vl_types.all;
entity RegResto_vlg_vec_tst is
end RegResto_vlg_vec_tst;
