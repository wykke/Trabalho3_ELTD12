library verilog;
use verilog.vl_types.all;
entity AntiLoopM_vlg_vec_tst is
end AntiLoopM_vlg_vec_tst;
