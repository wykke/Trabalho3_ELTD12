library verilog;
use verilog.vl_types.all;
entity SISTEMA_FINAL_vlg_vec_tst is
end SISTEMA_FINAL_vlg_vec_tst;
