library verilog;
use verilog.vl_types.all;
entity AntiLoopD_vlg_vec_tst is
end AntiLoopD_vlg_vec_tst;
