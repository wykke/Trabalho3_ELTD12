library verilog;
use verilog.vl_types.all;
entity regA_vlg_vec_tst is
end regA_vlg_vec_tst;
