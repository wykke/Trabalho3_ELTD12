library verilog;
use verilog.vl_types.all;
entity regC_vlg_vec_tst is
end regC_vlg_vec_tst;
