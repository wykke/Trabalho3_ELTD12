library verilog;
use verilog.vl_types.all;
entity Sistema_TB is
end Sistema_TB;
