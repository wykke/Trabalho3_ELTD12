library verilog;
use verilog.vl_types.all;
entity AntiLoop_vlg_vec_tst is
end AntiLoop_vlg_vec_tst;
